--=============================================================================
--Library Declarations:
--=============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;
library UNISIM;
use UNISIM.VComponents.all;
--=============================================================================
--Entity Declaration:
--=============================================================================
entity {component_name}_tb is
end entity;
--=============================================================================
--Architecture
--=============================================================================
architecture testbench of {component_name}_tb is
--=============================================================================
--Component Declaration
--=============================================================================
component {component_name} is
    Generic (
    {generics}
    );
    Port ( 
    {ports}
    );
end component;
--=============================================================================
--Signals
--=============================================================================
{internal_signals}
begin
--=============================================================================
--Port Map
--=============================================================================
uut: {component_name} 
	port map(		
  {port_connections}
  );
--=============================================================================
--clk_100MHz generation 
--=============================================================================
clkgen_proc: process
begin
{clk_gen}
end process clkgen_proc;
--=============================================================================
--Stimulus Process
--=============================================================================
stim_proc: process
begin				
{stim_proc}
wait;
end process stim_proc;
end testbench;
